`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/12/12 11:38:29
// Design Name: 
// Module Name: Mem_reg_WB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Mem_reg_WB(
    input wire clk_MemWB,
    input wire rst_MemWB,
    input wire en_MemWB,
    input wire valid_in_MemWB,//new
    input wire [31:0] PC4_in_MemWB,
    input wire [4:0] Rd_addr_MemWB,
    input wire [31:0] ALU_in_MemWB,
    input wire [31:0] DMem_data_MemWB,
    input wire [1:0] MemtoReg_in_MemWB,
    input wire RegWrite_in_MemWB,
    input wire [31:0] pc_in_MemWB,
    input wire [31:0] inst_in_MemWB,///
    output reg [31:0] PC4_out_MemWB,
    output reg [4:0] Rd_addr_out_MemWB,
    output reg [31:0] ALU_out_MemWB,
    output reg [31:0] DMem_data_out_MemWB,
    output reg [1:0] MemtoReg_out_MemWB,
    output reg RegWrite_out_MemWB,
    output reg [31:0] pc_out_MemWB,
    output reg [31:0] inst_out_MemWB,
    output reg valid_out_MemWB//new
    );
    
    always @ (posedge clk_MemWB or posedge rst_MemWB) begin
        if(en_MemWB == 1'b1) begin
            if(rst_MemWB == 1'b1) begin
                PC4_out_MemWB <= 32'b0;
                Rd_addr_out_MemWB <= 5'b0;
                ALU_out_MemWB <= 32'b0;
                DMem_data_out_MemWB <= 32'b0;
                MemtoReg_out_MemWB <= 2'b0;
                RegWrite_out_MemWB <= 1'b0;
                pc_out_MemWB <= 32'b0;
                inst_out_MemWB <= 32'b0;
                valid_out_MemWB <= valid_in_MemWB;
            end else begin
                PC4_out_MemWB <= PC4_in_MemWB;
                Rd_addr_out_MemWB <= Rd_addr_MemWB;
                ALU_out_MemWB <= ALU_in_MemWB;
                DMem_data_out_MemWB <= DMem_data_MemWB;
                MemtoReg_out_MemWB <= MemtoReg_in_MemWB;
                RegWrite_out_MemWB <= RegWrite_in_MemWB;
                pc_out_MemWB <= pc_in_MemWB;
                inst_out_MemWB <= inst_in_MemWB;
                valid_out_MemWB <= valid_in_MemWB;
            end
        end
    end
endmodule
