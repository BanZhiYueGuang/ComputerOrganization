module ADC_32(
    input [31:0] A,
    input [31:0] B,
    input C0,
    output [32:0] O
);

    // �� C0=1 ʱִ�м�����C0=0 ʱִ�мӷ�
    wire [31:0] B_modified;

    assign B_modified = C0 ? ~B : B;  // ����ʱȡ��B
    assign O = {1'b0, A} + {1'b0, B_modified} + C0; // ִ�мӷ�����

endmodule